module and_gate(a,b,y);
input a,b;
output y;
and a1(y,a,b);
endmodule

